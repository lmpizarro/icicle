// Defines for EDU-FPGA
